module CODEC
(
    input clk,
    input rst_n,

    input out,
    input en,
    input samp,

    output AUD_ADCLRCK,
    output AUD_ADCDAT,
    output AUD_DACLRCK,
    output AUD_DACDAT,
    output AUD_XCK,
    output AUD_BCLK,
    output I2C_SCLK,
    output I2C_SDAT
);

endmodule