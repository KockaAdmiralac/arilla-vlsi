module morse_code_receive_rom
(
	input      [7:0] in,
	output reg [7:0] out
);

always @(*)
begin
	case(in)
		8'b010_00001: out = 8'h41;//A
		8'b100_01000: out = 8'h42;//B
		8'b100_01010: out = 8'h43;//C
		8'b011_00100: out = 8'h44;//D
		8'b001_00000: out = 8'h45;//E
		8'b100_00010: out = 8'h46;//F
		8'b011_00110: out = 8'h47;//G
		8'b100_00000: out = 8'h48;//H
		8'b010_00000: out = 8'h49;//I
		8'b100_00111: out = 8'h4A;//J
		8'b011_00101: out = 8'h4B;//K
		8'b100_00100: out = 8'h4C;//L
		8'b010_00011: out = 8'h4D;//M
		8'b010_00010: out = 8'h4E;//N
		8'b011_00111: out = 8'h4F;//O
		8'b100_00110: out = 8'h50;//P
		8'b100_01101: out = 8'h51;//Q
		8'b011_00010: out = 8'h52;//R
		8'b011_00000: out = 8'h53;//S
		8'b001_00001: out = 8'h54;//T
		8'b011_00001: out = 8'h55;//U
		8'b100_00001: out = 8'h56;//V
		8'b011_00011: out = 8'h57;//W
		8'b100_01001: out = 8'h58;//X
		8'b100_01011: out = 8'h59;//Y
		8'b100_01100: out = 8'h5A;//Z
		8'b101_11111: out = 8'h30;//0
		8'b101_01111: out = 8'h31;//1
		8'b101_00111: out = 8'h32;//2
		8'b101_00011: out = 8'h33;//3
		8'b101_00001: out = 8'h34;//4
		8'b101_00000: out = 8'h35;//5
		8'b101_10000: out = 8'h36;//6
		8'b101_11000: out = 8'h37;//7
		8'b101_11100: out = 8'h38;//8
		8'b101_11110: out = 8'h39;//9
		8'b110_00000: out = 8'h20;//' '
		8'b111_00000: out = 8'h03;//ETX
		default:      out = 8'h00;
	endcase
end

endmodule