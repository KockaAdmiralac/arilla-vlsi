module SRAM
(
    input [3:0] ByteEna,
    input clk,

    input RD,
    input WR,
    input [31:0] ADDR,
    inout [31:0] DATA
);

endmodule