module MC_ROM
(
	input [7:0] in,
	output reg [7:0] out
);
	always @(*)
	begin
		case (in)
			8'h41: out = 8'b010_00001;//A
			8'h42: out = 8'b100_01000;//B
			8'h43: out = 8'b100_01010;//C
			8'h44: out = 8'b011_00100;//D
			8'h45: out = 8'b001_00000;//E
			8'h46: out = 8'b100_00010;//F
			8'h47: out = 8'b011_00110;//G
			8'h48: out = 8'b100_00000;//H
			8'h49: out = 8'b010_00000;//I
			8'h4A: out = 8'b100_00111;//J
			8'h4B: out = 8'b011_00101;//K
			8'h4C: out = 8'b100_00100;//L
			8'h4D: out = 8'b010_00011;//M
			8'h4E: out = 8'b010_00010;//N
			8'h4F: out = 8'b011_00111;//O
			8'h50: out = 8'b100_00110;//P
			8'h51: out = 8'b100_01101;//Q
			8'h52: out = 8'b011_00010;//R
			8'h53: out = 8'b011_00000;//S
			8'h54: out = 8'b001_00001;//T
			8'h55: out = 8'b011_00001;//U
			8'h56: out = 8'b100_00001;//V
			8'h57: out = 8'b011_00011;//W
			8'h58: out = 8'b100_01001;//X
			8'h59: out = 8'b100_01011;//Y
			8'h5A: out = 8'b100_01100;//Z
			8'h30: out = 8'b101_11111;//0
			8'h31: out = 8'b101_01111;//1
			8'h32: out = 8'b101_00111;//2
			8'h33: out = 8'b101_00011;//3
			8'h34: out = 8'b101_00001;//4
			8'h35: out = 8'b101_00000;//5
			8'h36: out = 8'b101_10000;//6
			8'h37: out = 8'b101_11000;//7
			8'h38: out = 8'b101_11100;//8
			8'h39: out = 8'b101_11110;//9
			8'h20: out = 8'b110_00000;//' '
			8'h03: out = 8'b111_00000;//ETX
			default: out=8'b000_00000;
		endcase
	end
endmodule