module PS2_keyboard_controller 
(
    input K_CLK,
    input K_DATA,
    input clk,
    input rst_n,
    output [23:0] K_CD,
    output P_ERR,
    output F_ERR
);
    
endmodule